library verilog;
use verilog.vl_types.all;
entity sopc_min is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
end sopc_min;
